module bad_alu;
    logic a;

    assign b = a;   // Error: 'b' is not declared

endmodule
