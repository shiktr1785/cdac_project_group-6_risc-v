
`ifndef INSTR_MEM_PKG_SV
`define INSTR_MEM_PKG_SV

package instr_mem_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"
    `include "instr_mem_seq_item.sv"
    `include "instr_mem_sequence.sv"
    
endpackage: instr_mem_pkg

`endif