`ifndef __PARAMS_SVH
`define __PARAMS_SVH

parameter int DATA_WIDTH   = 32;
parameter int OPCODE_WIDTH = 4;

`endif
