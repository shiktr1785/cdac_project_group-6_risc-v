// Code your design here
module top(
		input bit clock,
		input reset_n
);
  
  // Internal Wires & Buses
  
  // Instruction Memory Interface
  logic [31:0] instr;
  logic        instr_valid;
  logic        next_instr;
  
  // Decoder
  logic [3:0]  opcode;
  logic [31:0] imme_data;
  logic        rd2_imme_sel;
  logic [14:0] rs1_rs2_rd;
  logic        rs_addr_valid;
  logic        rs_store;
  logic        rd_wr_en;
  
  // Mux Output
  logic [31:0] imme_rs;
  
  // Register File Data
  logic [31:0] rs_data;      
  logic [31:0] rs_data_mux;   
  logic        op_done;
  
  // ALU Interface 
  logic [31:0] alu_data_out;
  logic        alu_data_valid;
  
  logic final_wr_en;
  assign final_wr_en = rd_wr_en & alu_data_valid;
  
  logic        op_done_final;
  assign op_done_final = op_done;
  
  // rd2_imme_sel - 0 for imme, 1 for rs2
  assign w_imme_rs = (w_rd2_imme_sel) ? w_rs_data_mux : w_imme_data;
  
  // Module Instantiations
  
  // 1) Instruction Memory
  instr_mem_v1 #(
        .DEPTH(64)          
  ) i_inst_mem (
        .clk        (clk),
        .reset_n    (reset_n),
        .next_instr (next_instr),   // Input from Decoder
        .instr      (instr),        // Output to Decoder
        .instr_valid(instr_valid)   // Output to Decoder
    );
  
  // 2) Decoder
  decoder_v2 i_decoder (
        .clk            (clk),
        .reset_n        (reset_n),
        .instr          (instr),
        .instr_valid    (instr_valid),
    	// To RegFile's op_done
    	.op_done        (op_done_final),      
        
        .next_instr     (next_instr),
        .opcode         (opcode),
        .imme_data      (imme_data),
        .rd2_imme_sel   (rd2_imme_sel),
        .rs1_rs2_rd     (rs1_rs2_rd),
        .rs_addr_valid  (rs_addr_valid),
        .rs_store       (rs_store),
        .rd_wr_en       (rd_wr_en)
    );
  
  // 3) Reg File
  reg_file i_regfile (
        .clk            (clk),
        .reset_n        (reset_n),
    
        // Controls
        .rs_addr_valid  (rs_addr_valid),
        .rs1_rs2_rd     (rs1_rs2_rd),
        .rd_wr_en       (final_wr_en),
        .rs_store       (rs_store),
    
    	// For immediate store
        .imme_data      (imme_data), 
    
        // Write back data from ALU
        .alu_data_out   (alu_data_out), 
        
    	.rs_data        (rs_data),      // Connected to ALU 
        .rs_data_mux    (rs_data_mux),  // Connected to Mux 
        .op_done        (op_done)       // Connected to Decoder
    );
  
  // 4) ALU
 	alu i_alu (
   		.rs_data        (rs_data),     // Operand 1 -from RegFile
   		.imme_rs        (imme_rs),      // Operand 2 - from Mux
   		.opcode         (opcode),       // Control - from Decoder
   		.alu_data_out   (alu_data_out), // Result - to RegFile
        .alu_data_valid (alu_data_valid)// Status 
    );

endmodule

