module bad_alu;
    logic a = 1'b0;
    logic c;

    assign c = ~a;
endmodule
