`ifndef __PARAMS_SVH
`define __PARAMS_SVH

parameter ADDR_WIDTH = 15;
parameter BUS_WIDTH = 32;
parameter OPCODE_WIDTH = 4;
parameter DEPTH = 64;

`endif
