module bad_alu(input logic a, output logic c);

    assign c = ~a;
endmodule
