module bad_alu;

    logic a;

    assign b = a; // 'b' is not declared
    
endmodule