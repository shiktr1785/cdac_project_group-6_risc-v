/* verilator lint_off MULTITOP*/
`include "rtl/alu/alu.sv"
`include "rtl/instr_mem/instr_mem_v1.sv"
`include "rtl/regfile/regfile.sv"
`include "rtl/decoder/decoder_v2.sv"

/*verilator lint_on MULTITOP*/

