`ifndef __PARAMS_SVH
`define __PARAMS_SVH

parameter ADDR_WIDTH = 5;
parameter BUS_WIDTH = 32;
parameter OPCODE_WIDTH = 11;

`endif
