/* verilator lint_off MULTITOP*/
`include "alu.sv"
`include "instr_mem_v2.sv"
`include "regfile.sv"
`include "decoder_v2.sv"

/*verilator lint_on MULTITOP*/

